`default_nettype none
`timescale 1ns / 1ps

module EsdkTestbild(
	clk
);

input clk;

endmodule;

